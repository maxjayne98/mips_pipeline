`timescale 1ns/1ns

module DataMem(input[31:0] Address, write_d, input clk, rst, MemRead, MemWrite, output logic[31:0] read_d);
	logic[31:0] DMem[511:0];
	assign read_d= DMem[Address];
	
	// logic[31:0] modified_address;
	
	always@ (posedge clk, posedge rst) begin 
		// modified_address <= Address >> 1;
		DMem[251] <= 32'b 00000000000000000000000000000001;
		DMem[252] <= 32'b 00000000000000000000000000000010;
		DMem[253] <= 32'b 00000000000000000000000000000011;
		DMem[254] <= 32'b 00000000000000000000000000000100;
		DMem[255] <= 32'b 00000000000000000000000000000101;
		DMem[256] <= 32'b 00000000000000000000000000000110;
		DMem[257] <= 32'b 00000000000000000000000000000111;
		DMem[258] <= 32'b 00000000000000000000000000001000;
		DMem[259] <= 32'b 00000000000000000000000000001001;
		DMem[260] <= 32'b 00000000000000000000000000001010;

		DMem[261] <= 32'b 00000000000000000000000000001011;
		DMem[262] <= 32'b 00000000000000000000000000001100;
		DMem[263] <= 32'b 00000000000000000000000000001101;
		DMem[264] <= 32'b 00000000000000000000000000001110;
		DMem[265] <= 32'b 00000000000000000000000000001111;
		DMem[266] <= 32'b 00000000000000000000000000010000;
		DMem[267] <= 32'b 00000000000000000000000000010001;
		DMem[268] <= 32'b 00000000000000000000000000010010;
		DMem[269] <= 32'b 00000000000000000000000000010011;
		DMem[270] <= 32'b 00000000000000000000000000010100;
		// if (rst) begin 
		// 	integer i;
		// 	for(i=0; i<512; i=i+1)
		// 		DMem[i] <= 32'b0;
		// end
		if(MemWrite)
			DMem[Address] <= write_d;
	end	
endmodule 